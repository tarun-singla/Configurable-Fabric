//Test Bench
module FPGA_TB_1();
  
  reg [3:0] ra, rb;
  reg rci;
  wire [3:0] wsum;
  wire wco;
  
  reg [32:0] tb_mem [0:13];
  
//fpga(s0, s1, s2, s3, co, , , , , a0, a1, a2, a3, b0, b1, b2, b3, ci, , , , , )
  
  fpga fpga_inst(.o0(wsum[0]), .o1(wsum[1]), .o2(wsum[2]), .o3(wsum[3]), .o4(wco), .o5(), .o6(), .o7(), .o8(), .i0(ra[0]), .i1(ra[1]), .i2(ra[2]), .i3(ra[3]), .i4(rb[0]), .i5(rb[1]), .i6(rb[2]), .i7(rb[3]), .i8(rci), .i9(1'b0), .i10(1'b0), .i11(1'b0), .clear(1'b0), .clock(1'b0));
  
  initial $readmemh("configure1.mem", tb_mem);
  
  initial
    begin
      fpga_inst.select.mem = tb_mem[0];
      
      fpga_inst.lta_0.mem = tb_mem[1];
      fpga_inst.lta_1.mem = tb_mem[1];
      fpga_inst.lta_2.mem = tb_mem[1];
      fpga_inst.lta_3.mem = tb_mem[1];
      fpga_inst.lta_4.mem = tb_mem[1];
      fpga_inst.lta_5.mem = tb_mem[1];
      fpga_inst.lta_6.mem = tb_mem[1];
      fpga_inst.lta_7.mem = tb_mem[1];
      
      fpga_inst.sb0a.configure = tb_mem[2][15:0];
      fpga_inst.sb1a.configure = tb_mem[2][15:0];
      fpga_inst.sb2a.configure = tb_mem[2][15:0];
      fpga_inst.sb3a.configure = tb_mem[2][15:0];
      fpga_inst.sb4a.configure = tb_mem[2][15:0];
      fpga_inst.sb5a.configure = tb_mem[2][15:0];
      fpga_inst.sb6a.configure = tb_mem[2][15:0];
      fpga_inst.sb7a.configure = tb_mem[2][15:0];
      
      fpga_inst.sb0b.configure = tb_mem[2][15:0];
      fpga_inst.sb1b.configure = tb_mem[2][15:0];
      fpga_inst.sb2b.configure = tb_mem[2][15:0];
      fpga_inst.sb3b.configure = tb_mem[2][15:0];
      fpga_inst.sb4b.configure = tb_mem[2][15:0];
      fpga_inst.sb5b.configure = tb_mem[2][15:0];
      fpga_inst.sb6b.configure = tb_mem[2][15:0];
      fpga_inst.sb7b.configure = tb_mem[2][15:0];
      
      fpga_inst.sb0c.configure = tb_mem[2][15:0];
      fpga_inst.sb1c.configure = tb_mem[2][15:0];
      fpga_inst.sb2c.configure = tb_mem[2][15:0];
      fpga_inst.sb3c.configure = tb_mem[2][15:0];
      fpga_inst.sb4c.configure = tb_mem[2][15:0];
      fpga_inst.sb5c.configure = tb_mem[2][15:0];
      fpga_inst.sb6c.configure = tb_mem[2][15:0];
      fpga_inst.sb7c.configure = tb_mem[2][15:0];
      
      fpga_inst.sb0d.configure = tb_mem[3][15:0];
      fpga_inst.sb1d.configure = tb_mem[3][15:0];
      fpga_inst.sb2d.configure = tb_mem[3][15:0];
      fpga_inst.sb3d.configure = tb_mem[3][15:0];
      fpga_inst.sb4d.configure = tb_mem[3][15:0];
      fpga_inst.sb5d.configure = tb_mem[3][15:0];
      fpga_inst.sb6d.configure = tb_mem[3][15:0];
      fpga_inst.sb7d.configure = tb_mem[3][15:0];
      
      fpga_inst.lt_0.mem = tb_mem[4];
      fpga_inst.lt_1.mem = tb_mem[5];
      fpga_inst.lt_2.mem = tb_mem[6];
      fpga_inst.lt_3.mem = tb_mem[7];
      fpga_inst.lt_4.mem = tb_mem[8];
      fpga_inst.lt_5.mem = tb_mem[9];
      fpga_inst.lt_6.mem = tb_mem[10];
      fpga_inst.lt_7.mem = tb_mem[11];
      
      fpga_inst.sb0e.configure = tb_mem[12][15:0];
      fpga_inst.sb5e.configure = tb_mem[12][15:0];
      fpga_inst.sb6e.configure = tb_mem[12][15:0];
      fpga_inst.sb7e.configure = tb_mem[12][15:0];
      fpga_inst.sb8e.configure = tb_mem[12][15:0];
      
      fpga_inst.sb1e.configure = tb_mem[13][15:0];
      fpga_inst.sb2e.configure = tb_mem[13][15:0];
      fpga_inst.sb3e.configure = tb_mem[13][15:0];
      fpga_inst.sb4e.configure = tb_mem[13][15:0];
      
      ra = 4'b000; rb = 4'b0000; rci = 1'b0;
      #20
      $display("%b %b", wsum, wco);
      
      ra = 4'b1111; rb = 4'b1111; rci = 1'b1;
      #20
      $display("%b %b", wsum, wco);
      
      ra = 4'b0011; rb = 4'b0101; rci = 1'b0;
      #20
      $display("%b %b", wsum, wco);
      
      ra = 4'b1101; rb = 4'b0011; rci = 1'b1;
      #20
      $display("%b %b", wsum, wco);
      
    end
  
  initial
    begin
      $dumpfile("fpga.vcd");
      $dumpvars;
    end
  
endmodule